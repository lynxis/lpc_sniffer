module top #(parameter CLOCK_FREQ = 12000000, parameter BAUD_RATE = 115200)
(
	input [3:0] lpc_ad,
	input lpc_clock,
	input lpc_frame,
	input lpc_reset,
	input ext_clock,
	output uart_tx_pin,
	output lpc_clock_led,
	output lpc_frame_led,
	output lpc_reset_led,
	output valid_lpc_output_led,
	output overflow_led);

	/* power on reset */
	wire reset;

	/* buffering */
	wire [3:0] lpc_ad_buffered;
	wire lpc_clock_buffered;
	wire lpc_frame_buffered;
	wire lpc_reset_buffered;

	/* lpc */
	wire [3:0] dec_cyctype_dir;
	wire [31:0] dec_addr;
	wire [7:0] dec_data;

	/* bufferdomain*/
	wire [47:0] lpc_data;
	wire [47:0] write_data;
	wire lpc_data_enable;

	/* ring buffer */
	wire read_clock_enable;
	wire write_clock_enable;
	wire empty;
	wire overflow;

	/* mem2serial */
	wire [47:0] read_data;

	/* uart tx */
	wire uart_ready;
	wire [7:0] uart_data;
	wire uart_clock_enable;
	wire uart_clock;

	power_on_reset POR(
		.clock(ext_clock),
		.reset(reset));

	SB_GB AD0(
		.USER_SIGNAL_TO_GLOBAL_BUFFER(lpc_ad[0]),
		.GLOBAL_BUFFER_OUTPUT(lpc_ad_buffered[0]));
	SB_GB AD1(
		.USER_SIGNAL_TO_GLOBAL_BUFFER(lpc_ad[1]),
		.GLOBAL_BUFFER_OUTPUT(lpc_ad_buffered[1]));

	SB_GB AD2(
		.USER_SIGNAL_TO_GLOBAL_BUFFER(lpc_ad[2]),
		.GLOBAL_BUFFER_OUTPUT(lpc_ad_buffered[2]));

	SB_GB AD3(
		.USER_SIGNAL_TO_GLOBAL_BUFFER(lpc_ad[3]),
		.GLOBAL_BUFFER_OUTPUT(lpc_ad_buffered[3]));

	SB_GB CLOCK(
		.USER_SIGNAL_TO_GLOBAL_BUFFER(lpc_clock),
		.GLOBAL_BUFFER_OUTPUT(lpc_clock_buffered));
	SB_GB RESET(
		.USER_SIGNAL_TO_GLOBAL_BUFFER(lpc_reset),
		.GLOBAL_BUFFER_OUTPUT(lpc_reset_buffered));
	SB_GB FRAME(
		.USER_SIGNAL_TO_GLOBAL_BUFFER(lpc_frame),
		.GLOBAL_BUFFER_OUTPUT(lpc_frame_buffered));


	lpc LPC(
		.lpc_ad(lpc_ad_buffered),
		.lpc_clock(lpc_clock_buffered),
		.lpc_frame(lpc_frame_buffered),
		.lpc_reset(lpc_reset_buffered),
		.reset(reset),
		.out_cyctype_dir(dec_cyctype_dir),
		.out_addr(dec_addr),
		.out_data(dec_data),
		.out_clock_enable(lpc_data_enable));

	bufferdomain #(.AW(48))
		BUFFERDOMAIN(
			.input_data(lpc_data),
			.input_enable(lpc_data_enable),
			.reset(reset),
			.clock(ext_clock),
			.output_data(write_data),
			.output_enable(write_clock_enable));

	assign lpc_data[47:16] = dec_addr;
	assign lpc_data[15:8] = dec_data;
	assign lpc_data[7:4] = 0;
	assign lpc_data[3:0] = dec_cyctype_dir;

	ringbuffer #(.AW(10), .DW(48))
		RINGBUFFER (
			.reset(reset),
			.clock(ext_clock),
			.write_clock_enable(write_clock_enable),
			.read_clock_enable(read_clock_enable),
			.read_data(read_data),
			.write_data(write_data),
			.empty(empty),
			.overflow(overflow));

	mem2serial MEM_SERIAL(
		.reset(reset),
		.clock(ext_clock),
		.read_empty(empty),
		.read_clock_enable(read_clock_enable),
		.read_data(read_data),
		.uart_clock_enable(uart_clock_enable),
		.uart_ready(uart_ready),
		.uart_data(uart_data));

	uart_tx #(.CLOCK_FREQ(CLOCK_FREQ), .BAUD_RATE(BAUD_RATE))
		SERIAL (
			.read_data(uart_data),
			.read_clock_enable(uart_clock_enable),
			.reset(reset),
			.ready(uart_ready),
			.tx(uart_tx_pin),
			.clock(ext_clock),
			.uart_clock(uart_clock));

	trigger_led TRIGGERLPC(
		.reset(reset),
		.clock(ext_clock),
		.led(valid_lpc_output_led),
		.trigger(lpc_data_enable));

	assign lpc_clock_led = lpc_clock_buffered;
	assign lpc_frame_led = ~lpc_frame_buffered;
	assign lpc_reset_led = 1;
	assign overflow_led = overflow;
endmodule
